module google_custom_search

fn test_search() {
}
