module main

fn main() {
	println('ok')
}
