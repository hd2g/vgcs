module google_custom_search

import google_custom_search.api
import google_custom_search.response
import google_custom_search.query

pub struct Client {
}

// pub fn (self Client) search() !Response
